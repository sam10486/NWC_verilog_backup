`include "../include/define.svh"
`include "R16_BU.sv"
`include "R16_IN_mux.sv"

module R16_top(
    input clk,
    input rst, 
    input [`D_width-1:0] x0 ,
    input [`D_width-1:0] x1 ,
    input [`D_width-1:0] x2 ,
    input [`D_width-1:0] x3 ,
    input [`D_width-1:0] x4 ,
    input [`D_width-1:0] x5 ,
    input [`D_width-1:0] x6 ,
    input [`D_width-1:0] x7 ,
    input [`D_width-1:0] x8 ,
    input [`D_width-1:0] x9 ,
    input [`D_width-1:0] x10,
    input [`D_width-1:0] x11,
    input [`D_width-1:0] x12,
    input [`D_width-1:0] x13,
    input [`D_width-1:0] x14,
    input [`D_width-1:0] x15,

    input [`D_width-1:0] twiddle_0,
    input [`D_width-1:0] twiddle_1,
    input [`D_width-1:0] twiddle_2,
    input [`D_width-1:0] twiddle_3,
    input [`D_width-1:0] twiddle_4,
    input [`D_width-1:0] twiddle_5,
    input [`D_width-1:0] twiddle_6,
    input [`D_width-1:0] twiddle_7,
    input [`D_width-1:0] twiddle_8,
    input [`D_width-1:0] twiddle_9,
    input [`D_width-1:0] twiddle_10,
    input [`D_width-1:0] twiddle_11,
    input [`D_width-1:0] twiddle_12,
    input [`D_width-1:0] twiddle_13,
    input [`D_width-1:0] twiddle_14,
    input [`D_width-1:0] twiddle_15,

    input [`D_width-1:0] modulus,
    input ntt_enable,

    input [`D_width-1:0] R16_MA0_idx,
    input [`D_width-1:0] R16_MA1_idx,
    input [`D_width-1:0] R16_MA2_idx,
    input [`D_width-1:0] R16_MA3_idx,
    input [`D_width-1:0] R16_MA4_idx,
    input [`D_width-1:0] R16_MA5_idx,
    input [`D_width-1:0] R16_MA6_idx,
    input [`D_width-1:0] R16_MA7_idx,
    input [`D_width-1:0] R16_MA8_idx,
    input [`D_width-1:0] R16_MA9_idx,
    input [`D_width-1:0] R16_MA10_idx,
    input [`D_width-1:0] R16_MA11_idx,
    input [`D_width-1:0] R16_MA12_idx,
    input [`D_width-1:0] R16_MA13_idx,
    input [`D_width-1:0] R16_MA14_idx,
    input [`D_width-1:0] R16_MA15_idx,

    input [`D_width-1:0] R16_BN0_idx,
    input [`D_width-1:0] R16_BN1_idx,
    input [`D_width-1:0] R16_BN2_idx,
    input [`D_width-1:0] R16_BN3_idx,
    input [`D_width-1:0] R16_BN4_idx,
    input [`D_width-1:0] R16_BN5_idx,
    input [`D_width-1:0] R16_BN6_idx,
    input [`D_width-1:0] R16_BN7_idx,
    input [`D_width-1:0] R16_BN8_idx,
    input [`D_width-1:0] R16_BN9_idx,
    input [`D_width-1:0] R16_BN10_idx,
    input [`D_width-1:0] R16_BN11_idx,
    input [`D_width-1:0] R16_BN12_idx,
    input [`D_width-1:0] R16_BN13_idx,
    input [`D_width-1:0] R16_BN14_idx,
    input [`D_width-1:0] R16_BN15_idx,
    
    //output
    output logic [`D_width-1:0] y0,
    output logic [`D_width-1:0] y1,
    output logic [`D_width-1:0] y2,
    output logic [`D_width-1:0] y3,
    output logic [`D_width-1:0] y4,
    output logic [`D_width-1:0] y5,
    output logic [`D_width-1:0] y6,
    output logic [`D_width-1:0] y7,
    output logic [`D_width-1:0] y8,
    output logic [`D_width-1:0] y9,
    output logic [`D_width-1:0] y10,
    output logic [`D_width-1:0] y11,
    output logic [`D_width-1:0] y12,
    output logic [`D_width-1:0] y13,
    output logic [`D_width-1:0] y14,
    output logic [`D_width-1:0] y15,

    output logic ntt_done,

    output logic [`D_width-1:0] R16_MA0_idx_out ,
    output logic [`D_width-1:0] R16_MA1_idx_out ,
    output logic [`D_width-1:0] R16_MA2_idx_out ,
    output logic [`D_width-1:0] R16_MA3_idx_out ,
    output logic [`D_width-1:0] R16_MA4_idx_out ,
    output logic [`D_width-1:0] R16_MA5_idx_out ,
    output logic [`D_width-1:0] R16_MA6_idx_out ,
    output logic [`D_width-1:0] R16_MA7_idx_out ,
    output logic [`D_width-1:0] R16_MA8_idx_out ,
    output logic [`D_width-1:0] R16_MA9_idx_out ,
    output logic [`D_width-1:0] R16_MA10_idx_out,
    output logic [`D_width-1:0] R16_MA11_idx_out,
    output logic [`D_width-1:0] R16_MA12_idx_out,
    output logic [`D_width-1:0] R16_MA13_idx_out,
    output logic [`D_width-1:0] R16_MA14_idx_out,
    output logic [`D_width-1:0] R16_MA15_idx_out,

    output logic [`D_width-1:0] R16_BN0_idx_out ,
    output logic [`D_width-1:0] R16_BN1_idx_out ,
    output logic [`D_width-1:0] R16_BN2_idx_out ,
    output logic [`D_width-1:0] R16_BN3_idx_out ,
    output logic [`D_width-1:0] R16_BN4_idx_out ,
    output logic [`D_width-1:0] R16_BN5_idx_out ,
    output logic [`D_width-1:0] R16_BN6_idx_out ,
    output logic [`D_width-1:0] R16_BN7_idx_out ,
    output logic [`D_width-1:0] R16_BN8_idx_out ,
    output logic [`D_width-1:0] R16_BN9_idx_out ,
    output logic [`D_width-1:0] R16_BN10_idx_out,
    output logic [`D_width-1:0] R16_BN11_idx_out,
    output logic [`D_width-1:0] R16_BN12_idx_out,
    output logic [`D_width-1:0] R16_BN13_idx_out,
    output logic [`D_width-1:0] R16_BN14_idx_out,
    output logic [`D_width-1:0] R16_BN15_idx_out
);




    R16_BU R16_BU(
        x0 ,
        x1 ,
        x2 ,
        x3 ,
        x4 ,
        x5 ,
        x6 ,
        x7 ,
        x8 ,
        x9 ,
        x10,
        x11,
        x12,
        x13,
        x14,
        x15,
    );

endmodule