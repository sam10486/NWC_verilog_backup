`include "../include/define.svh"
`include "../mem/SRAM_DP_512.sv"